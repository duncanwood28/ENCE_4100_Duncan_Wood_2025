module char2seg(
	input 		[7:0] char,
	output reg	[7:0] HEX0
);

	wire [7:0] w_char;

	assign w_char = ((char >= 8'd65) && (char <= 8'd90)) ? (char + 8'd32 ) : char;

	always @(*) begin
	
		HEX0 = 8'hFF;
		
		// ASCII Table Mapping
		case(w_char)
			// Numbers
			8'd48: HEX0 = 8'b01000000; // 0
			8'd49: HEX0 = 8'b01111001; // 1
			8'd50: HEX0 = 8'b00100100; // 2
			8'd51: HEX0 = 8'b00110000; // 3
			8'd52: HEX0 = 8'b00011001; // 4
			8'd53: HEX0 = 8'b00010010; // 5
			8'd54: HEX0 = 8'b00000010; // 6
			8'd55: HEX0 = 8'b01111000; // 7
			8'd56: HEX0 = 8'b00000000; // 8
			8'd57: HEX0 = 8'b00011000; // 9
			// Letters
			8'd97: HEX0 = 8'b10001000; // a
			8'd98: HEX0 = 8'b10000011; // b
			8'd99: HEX0 = 8'b11000110; // c
			8'd100: HEX0 = 8'b10100001; // d
			8'd101: HEX0 = 8'b10000110; // E
			8'd102: HEX0 = 8'b10001110; // F
			8'd103: HEX0 = 8'b11000010; // G
			8'd104: HEX0 = 8'b10001001; // H
			8'd105: HEX0 = 8'b11111001; // I
			8'd106: HEX0 = 8'b11110001; // J
			8'd107: HEX0 = 8'b10011100; // k?
			8'd108: HEX0 = 8'b11000111; // L
			8'd109: HEX0 = 8'b10011100; // M?
			8'd110: HEX0 = 8'b10101011; // n
			8'd111: HEX0 = 8'b10100011; // o
			8'd112: HEX0 = 8'b10001100; // p
			8'd113: HEX0 = 8'b10011000; // q
			8'd114: HEX0 = 8'b10101111; // r
			8'd115: HEX0 = 8'b10010010; // s
			8'd116: HEX0 = 8'b11111000; // t
			8'd117: HEX0 = 8'b11100011; // u
			8'd118: HEX0 = 8'b10011100; // v?
			8'd119: HEX0 = 8'b10011100; // w?
			8'd120: HEX0 = 8'b10011100; // x?
			8'd121: HEX0 = 8'b10011100; // y?
			8'd122: HEX0 = 8'b10100100; // z
		endcase
	end

endmodule
